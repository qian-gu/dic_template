package blinky_pkg;

  parameter CNT_DW = 4;

endpackage
