//=============================================================================
// Filename      : blinky_pkg.sv
// Author        : Qian Gu
// Email         : guqian110@gmail.com
// Created on    : 2022-08-01 10:20:27 PM
// Last Modified : 2022-08-01 10:40:12 PM
//
//=============================================================================
//! blinky package
/// Contains all common parameters, type definations, and functions.
package blinky_pkg;

  /// Counter width
  parameter CounterWidth = 4;

endpackage
